module top_module (
    output out);

    buf(out, 1'b0);
    
endmodule
